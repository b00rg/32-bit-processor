----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 31.10.2024 13:47:07
-- Design Name: 
-- Module Name: DP_FunctionalUnit_22336157 - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity DP_FunctionalUnit_22336157 is
    Port ( B, A : in STD_LOGIC_VECTOR(31 downto 0);
        FS : in STD_LOGIC_VECTOR(4 downto 0);
        C, N, Z, V : out STD_LOGIC; 
        F : out STD_LOGIC_VECTOR(31 downto 0));
end DP_FunctionalUnit_22336157;



architecture Behavioral of DP_FunctionalUnit_22336157 is

begin


end Behavioral;
