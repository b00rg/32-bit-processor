-- 4 to 16
